// ----------------------------------------------------------------------------
// 
// 
// ----------------------------------------------------------------------------
module uart_tx #(
  parameter CLKDIV = 128
)(
  input clk,
  input rst,
  input tx_start,
  output tx_pin,
  output tx_busy,
  input [7:0] txdata
);

// ----------------------------------------------------------------------------
reg [$clog2(CLKDIV-1):0] txcnt;

// ----------------------------------------------------------------------------
reg tx_busy_reg;
reg [3:0] bitcnt;
reg [9:0] txdata_latched;

// ----------------------------------------------------------------------------
//
// ----------------------------------------------------------------------------
always @(posedge clk) begin
  // --------------------------------------------------------------------------
  if(rst == 1) begin
    txcnt <= 0;
    bitcnt <= 0;
    tx_busy <= 0;
    tx_busy_reg <= 0;
    txdata_latched <= {10'b1};
  // --------------------------------------------------------------------------
  //
  // --------------------------------------------------------------------------
  end else if(!tx_busy_reg) begin
    if(tx_start == 1) begin
      bitcnt <= 9;      
      txcnt <= (CLKDIV-1);
      tx_busy_reg <= 1;
      txdata_latched <= {1'd1, txdata, 1'b0}; // 1b STOP + 8b DATA + 1b START
    end
    tx_busy <= 0;
  // --------------------------------------------------------------------------
  //
  // --------------------------------------------------------------------------
  end else if(txcnt) begin
    txcnt <= txcnt - 1;
    tx_busy <= 1;
  // --------------------------------------------------------------------------
  // 
  // --------------------------------------------------------------------------
  end else begin
    if(bitcnt) begin
      bitcnt <= bitcnt - 1;
    end else begin
      tx_busy_reg <= 0;       
    end        
    txcnt <= (CLKDIV-1);
    txdata_latched = {1'b1, txdata_latched[8:1]};
  end
end

// ----------------------------------------------------------------------------
assign tx_pin = txdata_latched[0];

endmodule
