// ----------------------------------------------------------------------------
// 
// 
// ----------------------------------------------------------------------------
module uart_tx #(
  parameter CLKDIV = 128
)(
  input clk,
  input rst,
  input tx_start,
  output tx_pin,
  output reg tx_busy,
  input [7:0] txdata
);

// ----------------------------------------------------------------------------
reg [$clog2(CLKDIV-1):0] txcnt;

// ----------------------------------------------------------------------------
reg txFlag;
reg [3:0] bitcnt;
reg [9:0] txdata_latched;

// ----------------------------------------------------------------------------
assign tx_busy = tx_start ^ txFlag;

// ----------------------------------------------------------------------------
//
// ----------------------------------------------------------------------------
always @(posedge clk) begin
  // --------------------------------------------------------------------------
  if(rst == 1) begin
    txcnt <= 0;
    bitcnt <= 0;
    txFlag <= 0;
    txdata_latched <= {10'b1};
  // --------------------------------------------------------------------------
  //
  // --------------------------------------------------------------------------
  end else if(!txFlag) begin
    if(tx_start == 1) begin
      txFlag <= 1;
      bitcnt <= 9;      
      txcnt <= (CLKDIV-1);
      txdata_latched <= {1'd1, txdata, 1'b0}; // 1b STOP + 8b DATA + 1b START
    end
  // --------------------------------------------------------------------------
  //
  // --------------------------------------------------------------------------
  end else if(txcnt) begin
    txcnt <= txcnt - 1;
  // --------------------------------------------------------------------------
  // 
  // --------------------------------------------------------------------------
  end else begin
    if(bitcnt) begin
      bitcnt <= bitcnt - 1;
      txcnt <= (CLKDIV-1);
      txdata_latched <= {1'b1, txdata_latched[9:1]};
    end else begin
      txFlag <= 0;  
    end        
  end
end

// ----------------------------------------------------------------------------
assign tx_pin = txdata_latched[0];

endmodule
